`timescale 1ns / 1ps

module program_counter (in, out);
    input [63:0] in;
    output [63:0] out;
    
    
endmodule
